--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;

--entity To_SSD is
--  Port ( SyncK : in STD_LOGIC; -- 1 KHz Clock
--         First_Digit : in STD_LOGIC_VECTOR ( 3 downto 0);
--         Second_Digit : in STD_LOGIC_VECTOR ( 3 downto 0);
--         Third_Digit : in STD_LOGIC_VECTOR ( 3 downto 0);
--         Segment : out STD_LOGIC_VECTOR ( 6 downto 0); -- SSD output
--         an : out STD_LOGIC_VECTOR ( 3 downto 0) -- anode output
--        );
--end To_SSD;

--architecture Behavioral of To_SSD is

--    SHARED VARIABLE int : INTEGER := 0;
--    SIGNAL temp : STD_LOGIC_VECTOR ( 3 downto 0) := "0000";
----    SIGNAL Segment : STD_LOGIC_VECTOR ( 6 downto 0) := "1111110";
--    SIGNAL anode : STD_LOGIC_VECTOR ( 3 downto 0) := "1110";
--begin
    
----    seg <= Segment;
    
--    PROCESS (SyncK)
--    BEGIN
--        if ( SyncK'event and SyncK = '1') then
--            if ( int = 2) then
--                temp <= Third_Digit;
--                an <= "1011";
--                int := 0;
--            elsif ( int = 1) then
--                temp <= Second_Digit;
--                an <= "1101";
--                int := int + 1;
--            elsif ( int = 0) then
--                temp <= First_Digit;
--                an <= "1110";
--                int := int + 1;
--            end if;
--        end if;
--    END PROCESS;
    
--    PROCESS ( temp)
--    BEGIN
--        if ( temp = "0000") then
--            Segment <=  "1111110"; -- 0
--        elsif  ( temp = "0001") then
--            Segment <=  "0110000"; -- 1
--        elsif  ( temp = "0010") then
--            Segment <=  "1101101"; -- 2
--        elsif  ( temp = "0011") then
--            Segment <=  "1111001"; -- 3
--        elsif  ( temp = "0100") then
--            Segment <=  "0110011"; -- 4
--        elsif  ( temp = "0101") then
--            Segment <=  "1011011"; -- 5
--        elsif  ( temp = "0110") then
--            Segment <=  "1011111"; -- 6
--        elsif  ( temp = "0111") then
--            Segment <=  "1110000"; -- 7
--        elsif  ( temp = "1000") then
--            Segment <=  "1111111"; -- 8
--        elsif  ( temp = "1001") then
--            Segment <=  "1111011"; -- 9
--        end if;
--    END PROCESS;
--end Behavioral;