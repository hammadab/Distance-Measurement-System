---- 0 - NULL
---- 1 - 0
---- 2 - 1
---- 3 - 2
---- 4 - 3
---- 5 - 4
---- 6 - 5
---- 7 - 6
---- 8 - 7
---- 9 - 8
---- 10 - 9
---- 11 - =
---- 12 - A
---- 13 - B
---- 14 - C
---- 15 - D
---- 16 - E
---- 17 - F
---- 18 - G
---- 19 - H
---- 20 - I
---- 21 - J
---- 22 - K
---- 23 - L
---- 24 - M
---- 25 - N
---- 26 - O
---- 27 - P
---- 28 - Q
---- 29 - R
---- 30 - S
---- 31 - T
---- 32 - U
---- 33 - V
---- 34 - W
---- 35 - X
---- 36 - Y
---- 36 - Z

---- Block dimension = 8 x 16

--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;

--entity Fonts is
--  Port (    Char : in CHARACTER;
--            Char_0, Char_1, Char_2, Char_3, Char_4, Char_5, Char_6, Char_7, Char_8, Char_9, 
--            Char_a, Char_b, Char_c, Char_d, Char_e, Char_f : out STD_LOGIC_VECTOR ( 7 downto 0)
--        );
--end Fonts;

--architecture Behavioral of Fonts is
--    TYPE Char_Code is array ( 15 downto 0) of STD_LOGIC_VECTOR ( 7 downto 0);
--    TYPE Characters is array ( 37 downto 0) of Char_Code;
--    SIGNAL ROM : Characters := (   -- 2^11-by-8
--            -- NUL: code x00
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00000000", -- 2
--            "00000000", -- 3
--            "00000000", -- 4
--            "00000000", -- 5
--            "00000000", -- 6
--            "00000000", -- 7
--            "00000000", -- 8
--            "00000000", -- 9
--            "00000000", -- a
--            "00000000", -- b
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
----            -- EOT: code x04
----            ("00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00010000", -- 4    *
----            "00111000", -- 5   ***
----            "01111100", -- 6  *****
----            "11111110", -- 7 *******
----            "01111100", -- 8  *****
----            "00111000", -- 9   ***
----            "00010000", -- a    *
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- BEL: code x07
----            ("00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00000000", -- 5
----            "00011000", -- 6    **
----            "00111100", -- 7   ****
----            "00111100", -- 8   ****
----            "00011000", -- 9    **
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x0f
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00011000", -- 3    **
----            "00011000", -- 4    **
----            "11011011", -- 5 ** ** **
----            "00111100", -- 6   ****
----            "11100111", -- 7 ***  ***
----            "00111100", -- 8   ****
----            "11011011", -- 9 ** ** **
----            "00011000", -- a    **
----            "00011000", -- b    **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x16
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "11111110", -- 8 *******
----            "11111110", -- 9 *******
----            "11111110", -- a *******
----            "11111110", -- b *******
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x1a
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00011000", -- 5    **
----            "00001100", -- 6     **
----            "11111110", -- 7 *******
----            "00001100", -- 8     **
----            "00011000", -- 9    **
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x1b
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00110000", -- 5   **
----            "01100000", -- 6  **
----            "11111110", -- 7 *******
----            "01100000", -- 8  **
----            "00110000", -- 9   **
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x21
----            "00000000", -- 0
----            "00000000", -- 1
----            "00011000", -- 2    **
----            "00111100", -- 3   ****
----            "00111100", -- 4   ****
----            "00111100", -- 5   ****
----            "00011000", -- 6    **
----            "00011000", -- 7    **
----            "00011000", -- 8    **
----            "00000000", -- 9
----            "00011000", -- a    **
----            "00011000", -- b    **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x22
----            "00000000", -- 0
----            "01100110", -- 1  **  **
----            "01100110", -- 2  **  **
----            "01100110", -- 3  **  **
----            "00100100", -- 4   *  *
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00000000", -- 9
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x23
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "01101100", -- 3  ** **
----            "01101100", -- 4  ** **
----            "11111110", -- 5 *******
----            "01101100", -- 6  ** **
----            "01101100", -- 7  ** **
----            "01101100", -- 8  ** **
----            "11111110", -- 9 *******
----            "01101100", -- a  ** **
----            "01101100", -- b  ** **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x25
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "11000010", -- 4 **    *
----            "11000110", -- 5 **   **
----            "00001100", -- 6     **
----            "00011000", -- 7    **
----            "00110000", -- 8   **
----            "01100000", -- 9  **
----            "11000110", -- a **   **
----            "10000110", -- b *    **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x26
----            "00000000", -- 0
----            "00000000", -- 1
----            "00111000", -- 2   ***
----            "01101100", -- 3  ** **
----            "01101100", -- 4  ** **
----            "00111000", -- 5   ***
----            "01110110", -- 6  *** **
----            "11011100", -- 7 ** ***
----            "11001100", -- 8 **  **
----            "11001100", -- 9 **  **
----            "11001100", -- a **  **
----            "01110110", -- b  *** **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x27
----            "00000000", -- 0
----            "00110000", -- 1   **
----            "00110000", -- 2   **
----            "00110000", -- 3   **
----            "01100000", -- 4  **
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00000000", -- 9
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x28
----            "00000000", -- 0
----            "00000000", -- 1
----            "00001100", -- 2     **
----            "00011000", -- 3    **
----            "00110000", -- 4   **
----            "00110000", -- 5   **
----            "00110000", -- 6   **
----            "00110000", -- 7   **
----            "00110000", -- 8   **
----            "00110000", -- 9   **
----            "00011000", -- a    **
----            "00001100", -- b     **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x29
----            "00000000", -- 0
----            "00000000", -- 1
----            "00110000", -- 2   **
----            "00011000", -- 3    **
----            "00001100", -- 4     **
----            "00001100", -- 5     **
----            "00001100", -- 6     **
----            "00001100", -- 7     **
----            "00001100", -- 8     **
----            "00001100", -- 9     **
----            "00011000", -- a    **
----            "00110000", -- b   **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x2a
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "01100110", -- 5  **  **
----            "00111100", -- 6   ****
----            "11111111", -- 7 ********
----            "00111100", -- 8   ****
----            "01100110", -- 9  **  **
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x2b
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00011000", -- 5    **
----            "00011000", -- 6    **
----            "01111110", -- 7  ******
----            "00011000", -- 8    **
----            "00011000", -- 9    **
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x2c
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00011000", -- 9    **
----            "00011000", -- a    **
----            "00011000", -- b    **
----            "00110000", -- c   **
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x2d
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00000000", -- 5
----            "00000000", -- 6
----            "01111110", -- 7  ******
----            "00000000", -- 8
----            "00000000", -- 9
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x2e
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00000000", -- 9
----            "00011000", -- a    **
----            "00011000", -- b    **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x2f
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000010", -- 4       *
----            "00000110", -- 5      **
----            "00001100", -- 6     **
----            "00011000", -- 7    **
----            "00110000", -- 8   **
----            "01100000", -- 9  **
----            "11000000", -- a **
----            "10000000", -- b *
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
--            -- 0: code x30
--            ("00000000", -- 0
--            "00000000", -- 1
--            "01111100", -- 2  *****
--            "11000110", -- 3 **   **
--            "11000110", -- 4 **   **
--            "11001110", -- 5 **  ***
--            "11011110", -- 6 ** ****
--            "11110110", -- 7 **** **
--            "11100110", -- 8 ***  **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "01111100", -- b  *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- 1: code x31
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00011000", -- 2
--            "00111000", -- 3
--            "01111000", -- 4    **
--            "00011000", -- 5   ***
--            "00011000", -- 6  ****
--            "00011000", -- 7    **
--            "00011000", -- 8    **
--            "00011000", -- 9    **
--            "00011000", -- a    **
--            "01111110", -- b    **
--            "00000000", -- c    **
--            "00000000", -- d  ******
--            "00000000", -- e
--            "00000000"), -- f
--            -- 2: code x32
--            ("00000000", -- 0
--            "00000000", -- 1
--            "01111100", -- 2  *****
--            "11000110", -- 3 **   **
--            "00000110", -- 4      **
--            "00001100", -- 5     **
--            "00011000", -- 6    **
--            "00110000", -- 7   **
--            "01100000", -- 8  **
--            "11000000", -- 9 **
--            "11010110", -- a ** * **
--            "11101110", -- b *** ***
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- 3: code x33
--            ("00000000", -- 0
--            "00000000", -- 1
--            "01111100", -- 2  *****
--            "11000110", -- 3 **   **
--            "00000110", -- 4      **
--            "00000110", -- 5      **
--            "00111100", -- 6   ****
--            "00000110", -- 7      **
--            "00000110", -- 8      **
--            "00000110", -- 9      **
--            "11000110", -- a **   **
--            "01111100", -- b  *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- 4: code x34
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00001100", -- 2     **
--            "00011100", -- 3    ***
--            "00111100", -- 4   ****
--            "01101100", -- 5  ** **
--            "11001100", -- 6 **  **
--            "11111110", -- 7 *******
--            "00001100", -- 8     **
--            "00001100", -- 9     **
--            "00001100", -- a     **
--            "00011110", -- b    ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x35
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111110", -- 2 *******
--            "11000000", -- 3 **
--            "11000000", -- 4 **
--            "11000000", -- 5 **
--            "11111100", -- 6 ******
--            "00000110", -- 7      **
--            "00000110", -- 8      **
--            "00000110", -- 9      **
--            "11000110", -- a **   **
--            "01111100", -- b  *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x36
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00111000", -- 2   ***
--            "01100000", -- 3  **
--            "11000000", -- 4 **
--            "11000000", -- 5 **
--            "11111100", -- 6 ******
--            "11000110", -- 7 **   **
--            "11000110", -- 8 **   **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "01111100", -- b  *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x37
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111110", -- 2 *******
--            "11000110", -- 3 **   **
--            "00000110", -- 4      **
--            "00000110", -- 5      **
--            "00001100", -- 6     **
--            "00011000", -- 7    **
--            "00110000", -- 8   **
--            "00110000", -- 9   **
--            "00110000", -- a   **
--            "00110000", -- b   **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x38
--            ("00000000", -- 0
--            "00000000", -- 1
--            "01111100", -- 2  *****
--            "11000110", -- 3 **   **
--            "11000110", -- 4 **   **
--            "11000110", -- 5 **   **
--            "01111100", -- 6  *****
--            "11000110", -- 7 **   **
--            "11000110", -- 8 **   **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "01111100", -- b  *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x39
--            ("00000000", -- 0
--            "00000000", -- 1
--            "01111100", -- 2  *****
--            "11000110", -- 3 **   **
--            "11000110", -- 4 **   **
--            "11000110", -- 5 **   **
--            "01111110", -- 6  ******
--            "00000110", -- 7      **
--            "00000110", -- 8      **
--            "00000110", -- 9      **
--            "00001100", -- a     **
--            "01111000", -- b  ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
----            -- code x3a
----            ("00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00011000", -- 4    **
----            "00011000", -- 5    **
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00011000", -- 9    **
----            "00011000", -- a    **
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x3b
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00011000", -- 4    **
----            "00011000", -- 5    **
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00011000", -- 9    **
----            "00011000", -- a    **
----            "00110000", -- b   **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x3c
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000110", -- 3      **
----            "00001100", -- 4     **
----            "00011000", -- 5    **
----            "00110000", -- 6   **
----            "01100000", -- 7  **
----            "00110000", -- 8   **
----            "00011000", -- 9    **
----            "00001100", -- a     **
----            "00000110", -- b      **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
--            -- code x3d
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00000000", -- 2
--            "00000000", -- 3
--            "00000000", -- 4
--            "01111110", -- 5  ******
--            "00000000", -- 6
--            "00000000", -- 7
--            "01111110", -- 8  ******
--            "00000000", -- 9
--            "00000000", -- a
--            "00000000", -- b
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
----            -- code x3e
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "01100000", -- 3  **
----            "00110000", -- 4   **
----            "00011000", -- 5    **
----            "00001100", -- 6     **
----            "00000110", -- 7      **
----            "00001100", -- 8     **
----            "00011000", -- 9    **
----            "00110000", -- a   **
----            "01100000", -- b  **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x3f
----            "00000000", -- 0
----            "00000000", -- 1
----            "01111100", -- 2  *****
----            "11000110", -- 3 **   **
----            "11000110", -- 4 **   **
----            "00001100", -- 5     **
----            "00011000", -- 6    **
----            "00011000", -- 7    **
----            "00011000", -- 8    **
----            "00000000", -- 9
----            "00011000", -- a    **
----            "00011000", -- b    **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
--            -- A: code x41
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00010000", -- 2    *
--            "00111000", -- 3   ***
--            "01101100", -- 4  ** **
--            "11000110", -- 5 **   **
--            "11000110", -- 6 **   **
--            "11111110", -- 7 *******
--            "11000110", -- 8 **   **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "11000110", -- b **   **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            (-- B: code x42
--            "00000000", -- 0
--            "00000000", -- 1
--            "11111100", -- 2 ******
--            "01100110", -- 3  **  **
--            "01100110", -- 4  **  **
--            "01100110", -- 5  **  **
--            "01111100", -- 6  *****
--            "01100110", -- 7  **  **
--            "01100110", -- 8  **  **
--            "01100110", -- 9  **  **
--            "01100110", -- a  **  **
--            "11111100", -- b ******
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- C: code x43
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00111100", -- 2   ****
--            "01100110", -- 3  **  **
--            "11000010", -- 4 **    *
--            "11000000", -- 5 **
--            "11000000", -- 6 **
--            "11000000", -- 7 **
--            "11000000", -- 8 **
--            "11000010", -- 9 **    *
--            "01100110", -- a  **  **
--            "00111100", -- b   ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- D: code x44
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111000", -- 2 *****
--            "01101100", -- 3  ** **
--            "01100110", -- 4  **  **
--            "01100110", -- 5  **  **
--            "01100110", -- 6  **  **
--            "01100110", -- 7  **  **
--            "01100110", -- 8  **  **
--            "01100110", -- 9  **  **
--            "01101100", -- a  ** **
--            "11111000", -- b *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x45
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111110", -- 2 *******
--            "01100110", -- 3  **  **
--            "01100010", -- 4  **   *
--            "01101000", -- 5  ** *
--            "01111000", -- 6  ****
--            "01101000", -- 7  ** *
--            "01100000", -- 8  **
--            "01100010", -- 9  **   *
--            "01100110", -- a  **  **
--            "11111110", -- b *******
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x46
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111110", -- 2 *******
--            "01100110", -- 3  **  **
--            "01100010", -- 4  **   *
--            "01101000", -- 5  ** *
--            "01111000", -- 6  ****
--            "01101000", -- 7  ** *
--            "01100000", -- 8  **
--            "01100000", -- 9  **
--            "01100000", -- a  **
--            "11110000", -- b ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x47
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00111100", -- 2   ****
--            "01100110", -- 3  **  **
--            "11000010", -- 4 **    *
--            "11000000", -- 5 **
--            "11000000", -- 6 **
--            "11011110", -- 7 ** ****
--            "11000110", -- 8 **   **
--            "11000110", -- 9 **   **
--            "01100110", -- a  **  **
--            "00111010", -- b   *** *
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- H: code x48
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11000110", -- 2 **   **
--            "11000110", -- 3 **   **
--            "11000110", -- 4 **   **
--            "11000110", -- 5 **   **
--            "11111110", -- 6 *******
--            "11000110", -- 7 **   **
--            "11000110", -- 8 **   **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "11000110", -- b **   **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- I: code x49
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00111100", -- 2   ****
--            "00011000", -- 3    **
--            "00011000", -- 4    **
--            "00011000", -- 5    **
--            "00011000", -- 6    **
--            "00011000", -- 7    **
--            "00011000", -- 8    **
--            "00011000", -- 9    **
--            "00011000", -- a    **
--            "00111100", -- b   ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- J: code x4a
--            ("00000000", -- 0
--            "00000000", -- 1
--            "00011110", -- 2    ****
--            "00001100", -- 3     **
--            "00001100", -- 4     **
--            "00001100", -- 5     **
--            "00001100", -- 6     **
--            "00001100", -- 7     **
--            "11001100", -- 8 **  **
--            "11001100", -- 9 **  **
--            "11001100", -- a **  **
--            "01111000", -- b  ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- K: code x4b
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11100110", -- 2 ***  **
--            "01100110", -- 3  **  **
--            "01100110", -- 4  **  **
--            "01101100", -- 5  ** **
--            "01111000", -- 6  ****
--            "01111000", -- 7  ****
--            "01101100", -- 8  ** **
--            "01100110", -- 9  **  **
--            "01100110", -- a  **  **
--            "11100110", -- b ***  **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- L: code x4c
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11110000", -- 2 ****
--            "01100000", -- 3  **
--            "01100000", -- 4  **
--            "01100000", -- 5  **
--            "01100000", -- 6  **
--            "01100000", -- 7  **
--            "01100000", -- 8  **
--            "01100010", -- 9  **   *
--            "01100110", -- a  **  **
--            "11111110", -- b *******
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- M: code x4d
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11000011", -- 2 **    **
--            "11100111", -- 3 ***  ***
--            "11111111", -- 4 ********
--            "11111111", -- 5 ********
--            "11011011", -- 6 ** ** **
--            "11000011", -- 7 **    **
--            "11000011", -- 8 **    **
--            "11000011", -- 9 **    **
--            "11000011", -- a **    **
--            "11000011", -- b **    **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- N: code x4e
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11000110", -- 2 **   **
--            "11100110", -- 3 ***  **
--            "11110110", -- 4 **** **
--            "11111110", -- 5 *******
--            "11011110", -- 6 ** ****
--            "11001110", -- 7 **  ***
--            "11000110", -- 8 **   **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "11000110", -- b **   **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- O: code x4f
--            ("00000000", -- 0
--            "00000000", -- 1
--            "01111100", -- 2  *****
--            "11000110", -- 3 **   **
--            "11000110", -- 4 **   **
--            "11000110", -- 5 **   **
--            "11000110", -- 6 **   **
--            "11000110", -- 7 **   **
--            "11000110", -- 8 **   **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "01111100", -- b  *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- P: code x50
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111100", -- 2 ******
--            "01100110", -- 3  **  **
--            "01100110", -- 4  **  **
--            "01100110", -- 5  **  **
--            "01111100", -- 6  *****
--            "01100000", -- 7  **
--            "01100000", -- 8  **
--            "01100000", -- 9  **
--            "01100000", -- a  **
--            "11110000", -- b ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- Q: code x510
--            ("00000000", -- 0
--            "00000000", -- 1
--            "01111100", -- 2  *****
--            "11000110", -- 3 **   **
--            "11000110", -- 4 **   **
--            "11000110", -- 5 **   **
--            "11000110", -- 6 **   **
--            "11000110", -- 7 **   **
--            "11000110", -- 8 **   **
--            "11010110", -- 9 ** * **
--            "11011110", -- a ** ****
--            "01111100", -- b  *****
--            "00001100", -- c     **
--            "00001110", -- d     ***
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x52
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111100", -- 2 ******
--            "01100110", -- 3  **  **
--            "01100110", -- 4  **  **
--            "01100110", -- 5  **  **
--            "01111100", -- 6  *****
--            "01101100", -- 7  ** **
--            "01100110", -- 8  **  **
--            "01100110", -- 9  **  **
--            "01100110", -- a  **  **
--            "11100110", -- b ***  **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x53
--            ("00000000", -- 0
--            "00000000", -- 1
--            "01111100", -- 2  *****
--            "11000110", -- 3 **   **
--            "11000110", -- 4 **   **
--            "01100000", -- 5  **
--            "00111000", -- 6   ***
--            "00001100", -- 7     **
--            "00000110", -- 8      **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "01111100", -- b  *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x54
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111111", -- 2 ********
--            "11011011", -- 3 ** ** **
--            "10011001", -- 4 *  **  *
--            "00011000", -- 5    **
--            "00011000", -- 6    **
--            "00011000", -- 7    **
--            "00011000", -- 8    **
--            "00011000", -- 9    **
--            "00011000", -- a    **
--            "00111100", -- b   ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x55
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11000110", -- 2 **   **
--            "11000110", -- 3 **   **
--            "11000110", -- 4 **   **
--            "11000110", -- 5 **   **
--            "11000110", -- 6 **   **
--            "11000110", -- 7 **   **
--            "11000110", -- 8 **   **
--            "11000110", -- 9 **   **
--            "11000110", -- a **   **
--            "01111100", -- b  *****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x56
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11000011", -- 2 **    **
--            "11000011", -- 3 **    **
--            "11000011", -- 4 **    **
--            "11000011", -- 5 **    **
--            "11000011", -- 6 **    **
--            "11000011", -- 7 **    **
--            "11000011", -- 8 **    **
--            "01100110", -- 9  **  **
--            "00111100", -- a   ****
--            "00011000", -- b    **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x57
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11000011", -- 2 **    **
--            "11000011", -- 3 **    **
--            "11000011", -- 4 **    **
--            "11000011", -- 5 **    **
--            "11000011", -- 6 **    **
--            "11011011", -- 7 ** ** **
--            "11011011", -- 8 ** ** **
--            "11111111", -- 9 ********
--            "01100110", -- a  **  **
--            "01100110", -- b  **  **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x58
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11000011", -- 2 **    **
--            "11000011", -- 3 **    **
--            "01100110", -- 4  **  **
--            "00111100", -- 5   ****
--            "00011000", -- 6    **
--            "00011000", -- 7    **
--            "00111100", -- 8   ****
--            "01100110", -- 9  **  **
--            "11000011", -- a **    **
--            "11000011", -- b **    **
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x59
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11000011", -- 2 **    **
--            "11000011", -- 3 **    **
--            "11000011", -- 4 **    **
--            "01100110", -- 5  **  **
--            "00111100", -- 6   ****
--            "00011000", -- 7    **
--            "00011000", -- 8    **
--            "00011000", -- 9    **
--            "00011000", -- a    **
--            "00111100", -- b   ****
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000"), -- f
--            -- code x5a
--            ("00000000", -- 0
--            "00000000", -- 1
--            "11111111", -- 2 ********
--            "11000011", -- 3 **    **
--            "10000110", -- 4 *    **
--            "00001100", -- 5     **
--            "00111000", -- 6   ***
--            "00111000", -- 7   ***
--            "01100000", -- 8  **
--            "11000001", -- 9 **     *
--            "11000011", -- a **    **
--            "11111111", -- b ********
--            "00000000", -- c
--            "00000000", -- d
--            "00000000", -- e
--            "00000000") -- f
----            -- code x5b
----            "00000000", -- 0
----            "00000000", -- 1
----            "00111100", -- 2   ****
----            "00110000", -- 3   **
----            "00110000", -- 4   **
----            "00110000", -- 5   **
----            "00110000", -- 6   **
----            "00110000", -- 7   **
----            "00110000", -- 8   **
----            "00110000", -- 9   **
----            "00110000", -- a   **
----            "00111100", -- b   ****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x5c
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "10000000", -- 3 *
----            "11000000", -- 4 **
----            "11100000", -- 5 ***
----            "01110000", -- 6  ***
----            "00111000", -- 7   ***
----            "00011100", -- 8    ***
----            "00001110", -- 9     ***
----            "00000110", -- a      **
----            "00000010", -- b       *
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x5d
----            "00000000", -- 0
----            "00000000", -- 1
----            "00111100", -- 2   ****
----            "00001100", -- 3     **
----            "00001100", -- 4     **
----            "00001100", -- 5     **
----            "00001100", -- 6     **
----            "00001100", -- 7     **
----            "00001100", -- 8     **
----            "00001100", -- 9     **
----            "00001100", -- a     **
----            "00111100", -- b   ****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x5e
----            "00010000", -- 0    *
----            "00111000", -- 1   ***
----            "01101100", -- 2  ** **
----            "11000110", -- 3 **   **
----            "00000000", -- 4
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00000000", -- 9
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x5f
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00000000", -- 9
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "11111111", -- d ********
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x60
----            "00110000", -- 0   **
----            "00110000", -- 1   **
----            "00011000", -- 2    **
----            "00000000", -- 3
----            "00000000", -- 4
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00000000", -- 9
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- a: code x61
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "01111000", -- 5  ****
----            "00001100", -- 6     **
----            "01111100", -- 7  *****
----            "11001100", -- 8 **  **
----            "11001100", -- 9 **  **
----            "11001100", -- a **  **
----            "01110110", -- b  *** **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- b: code x62
----            "00000000", -- 0
----            "00000000", -- 1
----            "11100000", -- 2  ***
----            "01100000", -- 3   **
----            "01100000", -- 4   **
----            "01111000", -- 5   ****
----            "01101100", -- 6   ** **
----            "01100110", -- 7   **  **
----            "01100110", -- 8   **  **
----            "01100110", -- 9   **  **
----            "01100110", -- a   **  **
----            "01111100", -- b   *****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- c: code x63
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "01111100", -- 5  *****
----            "11000110", -- 6 **   **
----            "11000000", -- 7 **
----            "11000000", -- 8 **
----            "11000000", -- 9 **
----            "11000110", -- a **   **
----            "01111100", -- b  *****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- d: code x64
----            "00000000", -- 0
----            "00000000", -- 1
----            "00011100", -- 2    ***
----            "00001100", -- 3     **
----            "00001100", -- 4     **
----            "00111100", -- 5   ****
----            "01101100", -- 6  ** **
----            "11001100", -- 7 **  **
----            "11001100", -- 8 **  **
----            "11001100", -- 9 **  **
----            "11001100", -- a **  **
----            "01110110", -- b  *** **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- e: code x65
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "01111100", -- 5  *****
----            "11000110", -- 6 **   **
----            "11111110", -- 7 *******
----            "11000000", -- 8 **
----            "11000000", -- 9 **
----            "11000110", -- a **   **
----            "01111100", -- b  *****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- f: code x66
----            "00000000", -- 0
----            "00000000", -- 1
----            "00111000", -- 2   ***
----            "01101100", -- 3  ** **
----            "01100100", -- 4  **  *
----            "01100000", -- 5  **
----            "11110000", -- 6 ****
----            "01100000", -- 7  **
----            "01100000", -- 8  **
----            "01100000", -- 9  **
----            "01100000", -- a  **
----            "11110000", -- b ****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- g: code x67
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "01110110", -- 5  *** **
----            "11001100", -- 6 **  **
----            "11001100", -- 7 **  **
----            "11001100", -- 8 **  **
----            "11001100", -- 9 **  **
----            "11001100", -- a **  **
----            "01111100", -- b  *****
----            "00001100", -- c     **
----            "11001100", -- d **  **
----            "01111000", -- e  ****
----            "00000000"), -- f
----            -- h: code x68
----            "00000000", -- 0
----            "00000000", -- 1
----            "11100000", -- 2 ***
----            "01100000", -- 3  **
----            "01100000", -- 4  **
----            "01101100", -- 5  ** **
----            "01110110", -- 6  *** **
----            "01100110", -- 7  **  **
----            "01100110", -- 8  **  **
----            "01100110", -- 9  **  **
----            "01100110", -- a  **  **
----            "11100110", -- b ***  **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- i: code x69
----            "00000000", -- 0
----            "00000000", -- 1
----            "00011000", -- 2    **
----            "00011000", -- 3    **
----            "00000000", -- 4
----            "00111000", -- 5   ***
----            "00011000", -- 6    **
----            "00011000", -- 7    **
----            "00011000", -- 8    **
----            "00011000", -- 9    **
----            "00011000", -- a    **
----            "00111100", -- b   ****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- j: code x6a
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000110", -- 2      **
----            "00000110", -- 3      **
----            "00000000", -- 4
----            "00001110", -- 5     ***
----            "00000110", -- 6      **
----            "00000110", -- 7      **
----            "00000110", -- 8      **
----            "00000110", -- 9      **
----            "00000110", -- a      **
----            "00000110", -- b      **
----            "01100110", -- c  **  **
----            "01100110", -- d  **  **
----            "00111100", -- e   ****
----            "00000000"), -- f
----            -- k: code x6b
----            "00000000", -- 0
----            "00000000", -- 1
----            "11100000", -- 2 ***
----            "01100000", -- 3  **
----            "01100000", -- 4  **
----            "01100110", -- 5  **  **
----            "01101100", -- 6  ** **
----            "01111000", -- 7  ****
----            "01111000", -- 8  ****
----            "01101100", -- 9  ** **
----            "01100110", -- a  **  **
----            "11100110", -- b ***  **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- l: code x6c
----            "00000000", -- 0
----            "00000000", -- 1
----            "00111000", -- 2   ***
----            "00011000", -- 3    **
----            "00011000", -- 4    **
----            "00011000", -- 5    **
----            "00011000", -- 6    **
----            "00011000", -- 7    **
----            "00011000", -- 8    **
----            "00011000", -- 9    **
----            "00011000", -- a    **
----            "00111100", -- b   ****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- m: code x6d
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11100110", -- 5 ***  **
----            "11111111", -- 6 ********
----            "11011011", -- 7 ** ** **
----            "11011011", -- 8 ** ** **
----            "11011011", -- 9 ** ** **
----            "11011011", -- a ** ** **
----            "11011011", -- b ** ** **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- n: code x6e
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11011100", -- 5 ** ***
----            "01100110", -- 6  **  **
----            "01100110", -- 7  **  **
----            "01100110", -- 8  **  **
----            "01100110", -- 9  **  **
----            "01100110", -- a  **  **
----            "01100110", -- b  **  **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- o: code x6f
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "01111100", -- 5  *****
----            "11000110", -- 6 **   **
----            "11000110", -- 7 **   **
----            "11000110", -- 8 **   **
----            "11000110", -- 9 **   **
----            "11000110", -- a **   **
----            "01111100", -- b  *****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x70
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11011100", -- 5 ** ***
----            "01100110", -- 6  **  **
----            "01100110", -- 7  **  **
----            "01100110", -- 8  **  **
----            "01100110", -- 9  **  **
----            "01100110", -- a  **  **
----            "01111100", -- b  *****
----            "01100000", -- c  **
----            "01100000", -- d  **
----            "11110000", -- e ****
----            "00000000"), -- f
----            -- code x71
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "01110110", -- 5  *** **
----            "11001100", -- 6 **  **
----            "11001100", -- 7 **  **
----            "11001100", -- 8 **  **
----            "11001100", -- 9 **  **
----            "11001100", -- a **  **
----            "01111100", -- b  *****
----            "00001100", -- c     **
----            "00001100", -- d     **
----            "00011110", -- e    ****
----            "00000000"), -- f
----            -- code x72
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11011100", -- 5 ** ***
----            "01110110", -- 6  *** **
----            "01100110", -- 7  **  **
----            "01100000", -- 8  **
----            "01100000", -- 9  **
----            "01100000", -- a  **
----            "11110000", -- b ****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x73
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "01111100", -- 5  *****
----            "11000110", -- 6 **   **
----            "01100000", -- 7  **
----            "00111000", -- 8   ***
----            "00001100", -- 9     **
----            "11000110", -- a **   **
----            "01111100", -- b  *****
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x74
----            "00000000", -- 0
----            "00000000", -- 1
----            "00010000", -- 2    *
----            "00110000", -- 3   **
----            "00110000", -- 4   **
----            "11111100", -- 5 ******
----            "00110000", -- 6   **
----            "00110000", -- 7   **
----            "00110000", -- 8   **
----            "00110000", -- 9   **
----            "00110110", -- a   ** **
----            "00011100", -- b    ***
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x75
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11001100", -- 5 **  **
----            "11001100", -- 6 **  **
----            "11001100", -- 7 **  **
----            "11001100", -- 8 **  **
----            "11001100", -- 9 **  **
----            "11001100", -- a **  **
----            "01110110", -- b  *** **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x76
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11000011", -- 5 **    **
----            "11000011", -- 6 **    **
----            "11000011", -- 7 **    **
----            "11000011", -- 8 **    **
----            "01100110", -- 9  **  **
----            "00111100", -- a   ****
----            "00011000", -- b    **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x77
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11000011", -- 5 **    **
----            "11000011", -- 6 **    **
----            "11000011", -- 7 **    **
----            "11011011", -- 8 ** ** **
----            "11011011", -- 9 ** ** **
----            "11111111", -- a ********
----            "01100110", -- b  **  **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x78
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11000011", -- 5 **    **
----            "01100110", -- 6  **  **
----            "00111100", -- 7   ****
----            "00011000", -- 8    **
----            "00111100", -- 9   ****
----            "01100110", -- a  **  **
----            "11000011", -- b **    **
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x79
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11000110", -- 5 **   **
----            "11000110", -- 6 **   **
----            "11000110", -- 7 **   **
----            "11000110", -- 8 **   **
----            "11000110", -- 9 **   **
----            "11000110", -- a **   **
----            "01111110", -- b  ******
----            "00000110", -- c      **
----            "00001100", -- d     **
----            "11111000", -- e *****
----            "00000000"), -- f
----            -- code x7a
----            "00000000", -- 0
----            "00000000", -- 1
----            "00000000", -- 2
----            "00000000", -- 3
----            "00000000", -- 4
----            "11111110", -- 5 *******
----            "11001100", -- 6 **  **
----            "00011000", -- 7    **
----            "00110000", -- 8   **
----            "01100000", -- 9  **
----            "11000110", -- a **   **
----            "11111110", -- b *******
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x7b
----            "00000000", -- 0
----            "00000000", -- 1
----            "00001110", -- 2     ***
----            "00011000", -- 3    **
----            "00011000", -- 4    **
----            "00011000", -- 5    **
----            "01110000", -- 6  ***
----            "00011000", -- 7    **
----            "00011000", -- 8    **
----            "00011000", -- 9    **
----            "00011000", -- a    **
----            "00001110", -- b     ***
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x7d
----            "00000000", -- 0
----            "00000000", -- 1
----            "01110000", -- 2  ***
----            "00011000", -- 3    **
----            "00011000", -- 4    **
----            "00011000", -- 5    **
----            "00001110", -- 6     ***
----            "00011000", -- 7    **
----            "00011000", -- 8    **
----            "00011000", -- 9    **
----            "00011000", -- a    **
----            "01110000", -- b  ***
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
----            -- code x7e
----            "00000000", -- 0
----            "00000000", -- 1
----            "01110110", -- 2  *** **
----            "11011100", -- 3 ** ***
----            "00000000", -- 4
----            "00000000", -- 5
----            "00000000", -- 6
----            "00000000", -- 7
----            "00000000", -- 8
----            "00000000", -- 9
----            "00000000", -- a
----            "00000000", -- b
----            "00000000", -- c
----            "00000000", -- d
----            "00000000", -- e
----            "00000000"), -- f
--        );
        
--    SHARED VARIABLE index : INTEGER := 0;
--begin
    
--    process ( Char)
--    begin
--        if ( Char = '0') then
--            index := 1;
--        elsif ( Char = '1') then
--            index := 2;
--        elsif ( Char = '2') then
--            index := 3;
--        elsif ( Char = '3') then
--            index := 4;
--        elsif ( Char = '4') then
--            index := 5;
--        elsif ( Char = '5') then
--            index := 6;
--        elsif ( Char = '6') then
--            index := 7;
--        elsif ( Char = '7') then
--            index := 8;
--        elsif ( Char = '8') then
--            index := 9;
--        elsif ( Char = '9') then
--            index := 10;
--        elsif ( Char = '=') then
--            index := 11;
--        elsif ( Char = 'A') then
--            index := 12;
--        elsif ( Char = 'B') then
--            index := 13;
--        elsif ( Char = 'C') then
--            index := 14;
--        elsif ( Char = 'D') then
--            index := 15;
--        elsif ( Char = 'E') then
--            index := 16;
--        elsif ( Char = 'F') then
--            index := 17;
--        elsif ( Char = 'G') then
--            index := 18;
--        elsif ( Char = 'H') then
--            index := 19;
--        elsif ( Char = 'I') then
--            index := 20;
--        elsif ( Char = 'J') then
--            index := 21;
--        elsif ( Char = 'K') then
--            index := 22;
--        elsif ( Char = 'L') then
--            index := 23;
--        elsif ( Char = 'M') then
--            index := 24;
--        elsif ( Char = 'N') then
--            index := 25;
--        elsif ( Char = 'O') then
--            index := 26;
--        elsif ( Char = 'P') then
--            index := 27;
--        elsif ( Char = 'Q') then
--            index := 28;
--        elsif ( Char = 'R') then
--            index := 29;
--        elsif ( Char = 'S') then
--            index := 30;
--        elsif ( Char = 'T') then
--            index := 31;
--        elsif ( Char = 'U') then
--            index := 32;
--        elsif ( Char = 'V') then
--            index := 33;
--        elsif ( Char = 'W') then
--            index := 34;
--        elsif ( Char = 'X') then
--            index := 35;
--        elsif ( Char = 'Y') then
--            index := 36;
--        elsif ( Char = 'Z') then
--            index := 37;
--        else
--            index := 0;
--        end if;
--    end process;
    
--    Char_0 <= ROM( index)(0);
--    Char_1 <= ROM( index)(1);
--    Char_2 <= ROM( index)(2);
--    Char_3 <= ROM( index)(3);
--    Char_4 <= ROM( index)(4);
--    Char_5 <= ROM( index)(5);
--    Char_6 <= ROM( index)(6);
--    Char_7 <= ROM( index)(7);
--    Char_8 <= ROM( index)(8);
--    Char_9 <= ROM( index)(9);
--    Char_A <= ROM( index)(10);
--    Char_B <= ROM( index)(11);
--    Char_C <= ROM( index)(12);
--    Char_D <= ROM( index)(13);
--    Char_E <= ROM( index)(14);
--    Char_F <= ROM( index)(15);
--end Behavioral;